*** SPICE deck for cell TwoInAND{lay} from library 2InputAND
*** Created on Sat May 11, 2024 19:40:29
*** Last revised on Sun Aug 18, 2024 22:18:39
*** Written on Sun Aug 18, 2024 22:18:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: TwoInAND{lay}
Mnmos@0 gnd A net@0 gnd NMOS L=1.2U W=12U AS=23.22P AD=117.54P PS=27.6U PD=99U
Mnmos@1 net@0 B net@2 gnd NMOS L=1.2U W=12U AS=49.02P AD=23.22P PS=47.8U PD=27.6U
Mnmos@4 gnd net@2 out gnd NMOS L=1.2U W=6U AS=46.44P AD=117.54P PS=45.6U PD=99U
Mpmos@0 vdd A net@2 vdd PMOS L=1.2U W=12U AS=49.02P AD=105.42P PS=47.8U PD=91.4U
Mpmos@1 net@2 B vdd vdd PMOS L=1.2U W=12U AS=105.42P AD=49.02P PS=91.4U PD=47.8U
Mpmos@4 vdd net@2 out vdd PMOS L=1.2U W=12U AS=46.44P AD=105.42P PS=45.6U PD=91.4U

* Spice Code nodes in cell cell 'TwoInAND{lay}'
vdd vdd 0 DC 5
va A 0 pwl 10n 0 20n 5 40n 5 50n 0 70n 0 80n 5 100n 5 110n 0 130n 0 140n 5 160n 5 170n 0 190n 0 200n 5
vb B 0 pwl 10n 0 40n 0 50n 5 100n 5 110n 0 160n 0 170n 5 200n 5
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=4ns trag v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rais=1 td=4ns trag v(out) val=4.5 rais=1
.tran 0 250ns
.include "C:\Electric\C5_models.txt"
.END
