*** SPICE deck for cell 4Bit_OR{sch} from library 4Bit_OR
*** Created on Sun Aug 18, 2024 01:06:03
*** Last revised on Sun Aug 18, 2024 20:53:20
*** Written on Sun Aug 18, 2024 20:56:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 4Bit_OR{sch}
Mnmos@0 net@4 A gnd gnd NMOS L=1.2U W=6U
Mnmos@1 net@4 B gnd gnd NMOS L=1.2U W=6U
Mnmos@2 gnd C net@4 gnd NMOS L=1.2U W=6U
Mnmos@3 gnd D net@4 gnd NMOS L=1.2U W=6U
Mnmos@4 OUT net@4 gnd gnd NMOS L=1.2U W=12U
Mpmos@0 vdd A net@0 vdd PMOS L=1.2U W=12U
Mpmos@1 net@0 B net@1 vdd PMOS L=1.2U W=12U
Mpmos@2 net@46 C net@1 vdd PMOS L=1.2U W=12U
Mpmos@3 net@4 D net@46 vdd PMOS L=1.2U W=12U
Mpmos@4 vdd net@4 OUT vdd PMOS L=1.2U W=12U

* Spice Code nodes in cell cell '4Bit_OR{sch}'
vdd vdd 0 DC 5 
va3 A 0 pwl 10n 0 15n 0 30n 0 31n 0 50n 0 51n 5 70n 5
va2 B 0 pwl 10n 0 15n 0 30n 0 31n 0 50n 0 51n 0 70n 0
cload out 0 400fF 
.measure tran tf trig v(out) val=0.5 fall=1 td=4ns targ v(out) val=4.5 fall=1 
.measure tran tr trig v(out) val=0.5 rais=1 td=4ns targ v(out) val=4.5 rais=1 
.tran 80n .include C:\Electric\C5_models.txt
.END
